//aes top
//include both aes_cipher_top and aes_inv_cipher_top


